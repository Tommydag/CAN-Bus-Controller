`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:59:33 05/17/2015 
// Design Name: 
// Module Name:    bit_timing 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module bit_timing(
    input rx,
    input rst,
    input clk,
	output sampled_rx,
    output baud_clk
    );

	if(posedge reset





endmodule
